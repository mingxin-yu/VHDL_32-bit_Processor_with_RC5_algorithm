library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
entity IMEM is
port (
 PC_Address: in std_logic_vector(31 downto 0);
 instruction: out  std_logic_vector(31 downto 0)
);
end IMEM;

architecture Behavioral of IMEM is
signal IMEM_buffer_address: std_logic_vector(30 downto 0);
 --type ROM_type is array (0 to 2505 ) of std_logic_vector(15 downto 0);
 type ROM_type is array (0 to 2557 ) of std_logic_vector(15 downto 0);
 --type ROM_type is array (0 to 771 ) of std_logic_vector(15 downto 0);
 constant rom_data: ROM_type:=(
 "0000000000000000","0000000000000000", -- Input
 "0001110000010111","0000000001000000",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000110101",
 "0001110000010111","0000000001000001",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000110100",
 "0001110000010111","0000000001000010",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000110111",
 "0001110000010111","0000000001000011",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000110110",
 "0001110000010111","0000000001000100",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000111001",
 "0001110000010111","0000000001000101",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000111000",
 "0001110000010111","0000000001000110",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000111011",
 "0001110000010111","0000000001000111",
 "0001011011110111","0000000000010000",
 "0010000000010111","0000000000111010",
 "1111110000000000","0000000000000000",
 "0000000000000000","0000000000000000", -- Encoding
 "0001110000000001","0000000000111010",
 "0001010000100001","0000000000010000",
 "0001110000010101","0000000000111011",
 "0000000000110101","0000100000000001",
 "0001110000000010","0000000000111000",
 "0001010001000010","0000000000010000",
 "0001110000010101","0000000000111001",
 "0000000001010101","0001000000000001",
 "0001110000000101","0000000000000000",
 "0001010010100101","0000000000010000",
 "0001110000010101","0000000000000001",
 "0000000010110101","0010100000000001",
 "0001110000000110","0000000000000010",
 "0001010011000110","0000000000010000",
 "0001110000010101","0000000000000011",
 "0000000011010101","0011000000000001",
 "0000000000100101","0000100000000001",
 "0000000001000110","0001000000000001",
 "0000010000000011","0000000000000100",
 "0000010000000100","0000000000000110",
 "0000010000010100","0000000000110100",
 "0001110001100101","0000000000000000",
 "0001010010100101","0000000000010000",
 "0001110001110101","0000000000000001",
 "0000000010110101","0010100000000001",
 "0001110010000110","0000000000000000",
 "0001010011000110","0000000000010000",
 "0001110010010101","0000000000000001",
 "0000000011010101","0011000000000001",
 "0000000000100001","0011100000001001",
 "0000000001000010","0100000000001001",
 "0000000000100010","0100100000001001",
 "0000000011101000","0101000000001001",
 "0000000101001001","0101100000001001",
 "0000010000001100","0000000000011111",
 "0000110001001101","0000000000011111",
 "0000010101101111","0000000000000000",
 "0000010000010000","0000000000000001",
 "0001011000010000","0000000000011111",
 "0000010000001110","0000000000011111",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000000111100101","0000100000000001",
 "0000000000100001","0011100000001001",
 "0000000000100010","0100100000001001",
 "0000000011101000","0101000000001001",
 "0000000101001001","0101100000001001",
 "0000110000101101","0000000000011111",
 "0000010101101111","0000000000000000",
 "0000010000010000","0000000000000001",
 "0001011000010000","0000000000011111",
 "0000010000001110","0000000000011111",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000000111100110","0001000000000001",
 "0000010001100011","0000000000000100",
 "0000010010000100","0000000000000100",
 "0010101010000011","0000000000000010",
 "0011000000000000","0000000001100000", -- Jump 96
 "1111110000000000","0000000000000000",
 "0000000000000000","0000000000000000", -- Decoding
 "0001110000000001","0000000000111010",
 "0001010000100001","0000000000010000",
 "0001110000010101","0000000000111011",
 "0000000000110101","0000100000000001",
 "0001110000000010","0000000000111000",
 "0001010001000010","0000000000010000",
 "0001110000010101","0000000000111001",
 "0000000001010101","0001000000000001",
 "0000010000000011","0000000000110000",
 "0000010000000100","0000000000110010",
 "0001110001100101","0000000000000000",
 "0001010010100101","0000000000010000",
 "0001110001110101","0000000000000001",
 "0000000010110101","0010100000000001",
 "0001110010000110","0000000000000000",
 "0001010011000110","0000000000010000",
 "0001110010010101","0000000000000001",
 "0000000011010101","0011000000000001",
 "0000000001000110","0011100000000011",
 "0000010000001000","0000000000011111",
 "0000000000101000","0100100000000101",
 "0000010000001010","0000000000100000",
 "0000000101001001","0101100000000011",
 "0000000101101000","0101100000000101",
 "0000010000001101","0000000000000001",
 "0001010110101101","0000000000011111",
 "0000010011101100","0000000000000000",
 "0000010000001111","0000000000011111",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000000110001100","1000000000001001",
 "0000000000100001","1000100000001001",
 "0000000110000001","1001000000001001",
 "0000001000010001","1001100000001001",
 "0000001001110010","1010000000001001",
 "0000011010000010","0000000000000000",
 "0000000000100101","0011100000000011",
 "0000000001001000","0100100000000101",
 "0000000101001001","0101100000000011",
 "0000000101101000","0101100000000101",
 "0000010011101100","0000000000000000",
 "0000010000001111","0000000000011111",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000100111101111","0000000000000001",
 "0010010101101111","0000000000001000",
 "0000000110001101","0111000000000101",
 "0001010110001100","0000000000000001",
 "0010100000001110","0000000000000010",
 "0000010110001100","0000000000000001",
 "0000000110001100","1000000000001001",
 "0000000001000010","1000100000001001",
 "0000000110000010","1001000000001001",
 "0000001000010001","1001100000001001",
 "0000001001110010","1010000000001001",
 "0000011010000001","0000000000000000",
 "0000100001100011","0000000000000100",
 "0000100010000100","0000000000000100",
 "0001110001100101","0000000000000000",
 "0001010010100101","0000000000010000",
 "0001110001110101","0000000000000001",
 "0000000010110101","0010100000000001",
 "0001110010000110","0000000000000000",
 "0001010011000110","0000000000010000",
 "0001110010010101","0000000000000001",
 "0000000011010101","0011000000000001",
 "0010100001100000","0000000000000010",
 "0011000000000000","0000001110110000", -- jump 892 + 52 = 944
 "0001110001100101","0000000000000000",
 "0001010010100101","0000000000010000",
 "0001110001110101","0000000000000001",
 "0000000010110101","0010100000000001",
 "0001110010000110","0000000000000000",
 "0001010011000110","0000000000010000",
 "0001110010010101","0000000000000001",
 "0000000011010101","0011000000000001",
 "0000000001000110","0001000000000011",
 "0000000000100101","0000100000000011",
 "1111110000000000","0000000000000000",
 "0000000000000000","0000000000000000", --Key Gen
 "0001110000000001","0000000000111100",
 "0001010000100001","0000000000010000",
 "0001110000010101","0000000000111101",
 "0000000000110101","0000100000000001",
 "0001110000000010","0000000000111110",
 "0001010001000010","0000000000010000",
 "0001110000010101","0000000000111111",
 "0000000001010101","0001000000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000000000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000000001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000000010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000000011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000000100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000000101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000000110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000000111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000001000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000001001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000001010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000001011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000001100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000001101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000001110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000001111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000010000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000010001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000010010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000010011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000010100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000010101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000010110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000010111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000011000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000011001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000011010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000011011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000011100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000011101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000011110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000011111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000100000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000100001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000100010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000100011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000100100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000100101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000100110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000100111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000101000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000101001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000101010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000101011",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000101100",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000101101",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000101110",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000101111",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000110000",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000110001",
 "0000000000100010","0000100000000001",
 "0000000000100000","1011000000000001",
 "0010000000010110","0000000000110010",
 "0001011011010110","0000000000010000",
 "0010000000010110","0000000000110011",
 "0000010000000011","0000000000000000",
 "0000010000000100","0000000000000000",
 "0000010000000101","0000000000000000",
 "0000010000000110","0000000000110100",
 "0000010000000111","0000000000000000",
 "0000010000010010","0000000000110100",
 "0000010000010011","0000000000111100",
 "0000010000010100","0000000001001110",
 "0001110010101000","0000000000000000",
 "0001010100001000","0000000000010000",
 "0001110010110101","0000000000000001",
 "0000000100010101","0100000000000001",
 "0000000001100100","0100100000000001",
 "0000000100001001","0100000000000001",
 "0000010100001111","0000000000000000",
 "0000010000010000","0000000000000001",
 "0001011000010000","0000000000011111",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000010111101000","0000000000000000",
 "0000000100000000","1011000000000001",
 "0010000010110110","0000000000000000",
 "0001011011010110","0000000000010000",
 "0010000010110110","0000000000000001",
 "0000010100000011","0000000000000000",
 "0000000001100100","0100100000000001",
 "0000110100101010","0000000000011111",
 "0001110011001011","0000000000000000",
 "0001010101101011","0000000000010000",
 "0001110011010101","0000000000000001",
 "0000000101110101","0101100000000001",
 "0000000101101001","0101100000000001",
 "0000010101001101","0000000000000000",
 "0000010101101111","0000000000000000",
 "0000010000010000","0000000000000001",
 "0001011000010000","0000000000011111",
 "0000010000001110","0000000000011111",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000100111001110","0000000000000001",
 "0010010110101110","0000000000001000",
 "0000000111110000","1000100000000101",
 "0001010111101111","0000000000000001",
 "0010100000010001","0000000000000010",
 "0000010111101111","0000000000000001",
 "0000010111101011","0000000000000000",
 "0000000101100000","1011000000000001",
 "0010000011010110","0000000000000000",
 "0001011011010110","0000000000010000",
 "0010000011010110","0000000000000001",
 "0000010101100100","0000000000000000",
 "0000010011100111","0000000000000001",
 "0000010010100101","0000000000000010",
 "0000010011000110","0000000000000010",
 "0010010010110010","0000000000000010",
 "0000100010100101","0000000000110100",
 "0010010011010011","0000000000000010",
 "0000100011000110","0000000000001000",
 "0010101010000111","0000000000000010",
 "0011000000000000","0000100000011110",    -- jump 2026 + 52 = 2078
 "1111110000000000","0000000000000000"
  );

begin
IMEM_buffer_address <= PC_Address(31 downto 1);
instruction <= rom_data(CONV_INTEGER(IMEM_buffer_address(30 downto 0) & '0'))&rom_data(CONV_INTEGER(IMEM_buffer_address(30 downto 0) & '1'));
end Behavioral;