library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY Left_Rotate IS
  PORT (a: in STD_LOGIC_VECTOR(31 DOWNTO 0);
	   b: in STD_LOGIC_VECTOR(31 DOWNTO 0);
 	   o: out STD_LOGIC_VECTOR(31 DOWNTO 0));
END Left_Rotate;

ARCHITECTURE rtl OF Left_Rotate IS
--signal temp: STD_LOGIC_VECTOR (5 DOWNTO 0);
BEGIN
WITH b(4 DOWNTO 0) SELECT
    O<=	a(30 DOWNTO 0) & '0' WHEN "00001",
	a(29 DOWNTO 0) & "00" WHEN "00010",
	a(28 DOWNTO 0) & "000" WHEN "00011",
	a(27 DOWNTO 0) & "0000" WHEN "00100",
	a(26 DOWNTO 0) & "00000" WHEN "00101",
	a(25 DOWNTO 0) & "000000" WHEN "00110",
	a(24 DOWNTO 0) & "0000000" WHEN "00111",
	a(23 DOWNTO 0) & "00000000" WHEN "01000",
	a(22 DOWNTO 0) & "000000000" WHEN "01001",
	a(21 DOWNTO 0) & "0000000000" WHEN "01010",
	a(20 DOWNTO 0) & "00000000000" WHEN "01011",
	a(19 DOWNTO 0) & "000000000000" WHEN "01100",
	a(18 DOWNTO 0) & "0000000000000" WHEN "01101",
	a(17 DOWNTO 0) & "00000000000000" WHEN "01110",
	a(16 DOWNTO 0) & "000000000000000" WHEN "01111",
	a(15 DOWNTO 0) & "0000000000000000" WHEN "10000",
    a(14 DOWNTO 0) & "00000000000000000" WHEN "10001",
    a(13 DOWNTO 0) & "000000000000000000" WHEN "10010",
    a(12 DOWNTO 0) & "0000000000000000000" WHEN "10011",
    a(11 DOWNTO 0) & "00000000000000000000" WHEN "10100",
    a(10 DOWNTO 0) & "000000000000000000000" WHEN "10101",
    a(9 DOWNTO 0) &  "0000000000000000000000" WHEN "10110",
    a(8 DOWNTO 0) &  "00000000000000000000000" WHEN "10111",
    a(7 DOWNTO 0) &  "000000000000000000000000" WHEN "11000",
    a(6 DOWNTO 0) &  "0000000000000000000000000" WHEN "11001",
    a(5 DOWNTO 0) &  "00000000000000000000000000" WHEN "11010",
    a(4 DOWNTO 0) &  "000000000000000000000000000" WHEN "11011",
    a(3 DOWNTO 0) &  "0000000000000000000000000000" WHEN "11100",
    a(2 DOWNTO 0) &  "00000000000000000000000000000" WHEN "11101",
    a(1 DOWNTO 0) &  "000000000000000000000000000000" WHEN "11110",
    a(0) &           "0000000000000000000000000000000" WHEN "11111",
                     "00000000000000000000000000000000" WHEN OTHERS;
END rtl;